module I2S_Transmitter(
  input         clock,
  input         reset,
  input  [31:0] io_Tx,
  output        io_Ready,
  output        io_LRCLK,
  output        io_BCLK,
  output        io_MCLK,
  output [15:0] io_DATA,
  output        io_bDATA,
  output [1:0]  io_State_o,
  output [7:0]  io_BitCntr,
  output        io_tick,
  input  [15:0] io_sw,
  output [15:0] io_CLKR
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  pll_MCLK_48K; // @[Hello.scala 47:19]
  wire  pll_MCLK_44K; // @[Hello.scala 47:19]
  wire  pll_locked; // @[Hello.scala 47:19]
  wire  pll_clk_in1; // @[Hello.scala 47:19]
  reg  current_state; // @[Hello.scala 56:30]
  reg [7:0] Bit_Counter; // @[Hello.scala 57:30]
  reg [7:0] ClkCntr; // @[Hello.scala 58:30]
  reg  Tckr; // @[Hello.scala 59:30]
  reg  BCLKTckr; // @[Hello.scala 60:30]
  reg  LRClkr; // @[Hello.scala 61:30]
  reg  bDATA; // @[Hello.scala 62:30]
  reg [15:0] DATA; // @[Hello.scala 63:30]
  reg [31:0] lutOut; // @[Hello.scala 64:30]
  reg [15:0] FRAME_NR; // @[Hello.scala 65:30]
  wire [7:0] _ClkCntr_T_1 = ClkCntr + 8'h1; // @[Hello.scala 81:24]
  wire  _T_1 = ClkCntr == 8'h40; // @[Hello.scala 85:19]
  wire  _T_2 = ClkCntr == 8'h20 | _T_1; // @[Hello.scala 84:28]
  wire  _GEN_0 = _T_2 ? ~BCLKTckr : BCLKTckr; // @[Hello.scala 85:29 87:22 60:30]
  wire [15:0] _FRAME_NR_T_1 = FRAME_NR + 16'h1; // @[Hello.scala 102:28]
  wire [5:0] _T_12 = 6'h20 - 6'h1; // @[Hello.scala 134:66]
  wire [7:0] _GEN_2046 = {{2'd0}, _T_12}; // @[Hello.scala 134:57]
  wire [15:0] _GEN_6 = 10'h1 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(16'sh0); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_7 = 10'h2 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_6); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_8 = 10'h3 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_7); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_9 = 10'h4 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_8); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_10 = 10'h5 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_9); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_11 = 10'h6 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_10); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_12 = 10'h7 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_11); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_13 = 10'h8 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_12); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_14 = 10'h9 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_13); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_15 = 10'ha == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_14); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_16 = 10'hb == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_15); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_17 = 10'hc == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_16); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_18 = 10'hd == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_17); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_19 = 10'he == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_18); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_20 = 10'hf == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_19); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_21 = 10'h10 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_20); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_22 = 10'h11 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_21); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_23 = 10'h12 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_22); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_24 = 10'h13 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_23); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_25 = 10'h14 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_24); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_26 = 10'h15 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_25); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_27 = 10'h16 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_26); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_28 = 10'h17 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_27); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_29 = 10'h18 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_28); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_30 = 10'h19 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_29); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_31 = 10'h1a == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_30); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_32 = 10'h1b == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_31); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_33 = 10'h1c == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_32); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_34 = 10'h1d == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_33); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_35 = 10'h1e == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_34); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_36 = 10'h1f == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_35); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_37 = 10'h20 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_36); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_38 = 10'h21 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_37); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_39 = 10'h22 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_38); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_40 = 10'h23 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_39); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_41 = 10'h24 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_40); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_42 = 10'h25 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_41); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_43 = 10'h26 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_42); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_44 = 10'h27 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_43); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_45 = 10'h28 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_44); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_46 = 10'h29 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_45); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_47 = 10'h2a == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_46); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_48 = 10'h2b == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_47); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_49 = 10'h2c == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_48); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_50 = 10'h2d == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_49); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_51 = 10'h2e == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_50); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_52 = 10'h2f == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_51); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_53 = 10'h30 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_52); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_54 = 10'h31 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_53); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_55 = 10'h32 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_54); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_56 = 10'h33 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_55); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_57 = 10'h34 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_56); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_58 = 10'h35 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_57); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_59 = 10'h36 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_58); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_60 = 10'h37 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_59); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_61 = 10'h38 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_60); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_62 = 10'h39 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_61); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_63 = 10'h3a == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_62); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_64 = 10'h3b == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_63); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_65 = 10'h3c == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_64); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_66 = 10'h3d == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_65); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_67 = 10'h3e == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_66); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_68 = 10'h3f == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_67); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_69 = 10'h40 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_68); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_70 = 10'h41 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_69); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_71 = 10'h42 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_70); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_72 = 10'h43 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_71); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_73 = 10'h44 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_72); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_74 = 10'h45 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_73); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_75 = 10'h46 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_74); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_76 = 10'h47 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_75); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_77 = 10'h48 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_76); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_78 = 10'h49 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_77); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_79 = 10'h4a == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_78); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_80 = 10'h4b == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_79); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_81 = 10'h4c == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_80); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_82 = 10'h4d == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_81); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_83 = 10'h4e == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_82); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_84 = 10'h4f == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_83); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_85 = 10'h50 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_84); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_86 = 10'h51 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_85); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_87 = 10'h52 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_86); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_88 = 10'h53 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_87); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_89 = 10'h54 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_88); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_90 = 10'h55 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_89); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_91 = 10'h56 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_90); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_92 = 10'h57 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_91); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_93 = 10'h58 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_92); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_94 = 10'h59 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_93); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_95 = 10'h5a == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_94); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_96 = 10'h5b == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_95); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_97 = 10'h5c == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_96); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_98 = 10'h5d == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_97); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_99 = 10'h5e == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_98); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_100 = 10'h5f == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_99); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_101 = 10'h60 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_100); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_102 = 10'h61 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_101); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_103 = 10'h62 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_102); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_104 = 10'h63 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_103); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_105 = 10'h64 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_104); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_106 = 10'h65 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_105); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_107 = 10'h66 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_106); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_108 = 10'h67 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_107); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_109 = 10'h68 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_108); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_110 = 10'h69 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_109); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_111 = 10'h6a == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_110); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_112 = 10'h6b == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_111); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_113 = 10'h6c == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_112); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_114 = 10'h6d == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_113); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_115 = 10'h6e == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_114); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_116 = 10'h6f == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_115); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_117 = 10'h70 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_116); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_118 = 10'h71 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_117); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_119 = 10'h72 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_118); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_120 = 10'h73 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_119); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_121 = 10'h74 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_120); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_122 = 10'h75 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_121); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_123 = 10'h76 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_122); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_124 = 10'h77 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_123); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_125 = 10'h78 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_124); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_126 = 10'h79 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_125); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_127 = 10'h7a == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_126); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_128 = 10'h7b == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_127); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_129 = 10'h7c == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_128); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_130 = 10'h7d == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_129); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_131 = 10'h7e == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_130); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_132 = 10'h7f == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_131); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_133 = 10'h80 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_132); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_134 = 10'h81 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_133); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_135 = 10'h82 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_134); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_136 = 10'h83 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_135); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_137 = 10'h84 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_136); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_138 = 10'h85 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_137); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_139 = 10'h86 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_138); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_140 = 10'h87 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_139); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_141 = 10'h88 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_140); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_142 = 10'h89 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_141); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_143 = 10'h8a == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_142); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_144 = 10'h8b == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_143); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_145 = 10'h8c == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_144); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_146 = 10'h8d == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_145); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_147 = 10'h8e == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_146); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_148 = 10'h8f == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_147); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_149 = 10'h90 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_148); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_150 = 10'h91 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_149); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_151 = 10'h92 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_150); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_152 = 10'h93 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_151); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_153 = 10'h94 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_152); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_154 = 10'h95 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_153); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_155 = 10'h96 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_154); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_156 = 10'h97 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_155); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_157 = 10'h98 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_156); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_158 = 10'h99 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_157); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_159 = 10'h9a == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_158); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_160 = 10'h9b == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_159); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_161 = 10'h9c == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_160); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_162 = 10'h9d == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_161); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_163 = 10'h9e == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_162); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_164 = 10'h9f == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_163); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_165 = 10'ha0 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_164); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_166 = 10'ha1 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_165); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_167 = 10'ha2 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_166); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_168 = 10'ha3 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_167); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_169 = 10'ha4 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_168); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_170 = 10'ha5 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_169); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_171 = 10'ha6 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_170); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_172 = 10'ha7 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_171); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_173 = 10'ha8 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_172); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_174 = 10'ha9 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_173); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_175 = 10'haa == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_174); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_176 = 10'hab == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_175); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_177 = 10'hac == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_176); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_178 = 10'had == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_177); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_179 = 10'hae == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_178); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_180 = 10'haf == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_179); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_181 = 10'hb0 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_180); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_182 = 10'hb1 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_181); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_183 = 10'hb2 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_182); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_184 = 10'hb3 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_183); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_185 = 10'hb4 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_184); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_186 = 10'hb5 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_185); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_187 = 10'hb6 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_186); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_188 = 10'hb7 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_187); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_189 = 10'hb8 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_188); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_190 = 10'hb9 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_189); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_191 = 10'hba == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_190); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_192 = 10'hbb == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_191); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_193 = 10'hbc == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_192); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_194 = 10'hbd == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_193); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_195 = 10'hbe == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_194); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_196 = 10'hbf == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_195); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_197 = 10'hc0 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_196); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_198 = 10'hc1 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_197); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_199 = 10'hc2 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_198); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_200 = 10'hc3 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_199); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_201 = 10'hc4 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_200); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_202 = 10'hc5 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_201); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_203 = 10'hc6 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_202); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_204 = 10'hc7 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_203); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_205 = 10'hc8 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_204); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_206 = 10'hc9 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_205); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_207 = 10'hca == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_206); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_208 = 10'hcb == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_207); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_209 = 10'hcc == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_208); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_210 = 10'hcd == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_209); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_211 = 10'hce == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_210); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_212 = 10'hcf == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_211); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_213 = 10'hd0 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_212); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_214 = 10'hd1 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_213); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_215 = 10'hd2 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_214); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_216 = 10'hd3 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_215); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_217 = 10'hd4 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_216); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_218 = 10'hd5 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_217); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_219 = 10'hd6 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_218); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_220 = 10'hd7 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_219); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_221 = 10'hd8 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_220); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_222 = 10'hd9 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_221); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_223 = 10'hda == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_222); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_224 = 10'hdb == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_223); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_225 = 10'hdc == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_224); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_226 = 10'hdd == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_225); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_227 = 10'hde == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_226); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_228 = 10'hdf == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_227); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_229 = 10'he0 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_228); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_230 = 10'he1 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_229); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_231 = 10'he2 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_230); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_232 = 10'he3 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_231); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_233 = 10'he4 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_232); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_234 = 10'he5 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_233); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_235 = 10'he6 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_234); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_236 = 10'he7 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_235); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_237 = 10'he8 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_236); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_238 = 10'he9 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_237); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_239 = 10'hea == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_238); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_240 = 10'heb == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_239); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_241 = 10'hec == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_240); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_242 = 10'hed == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_241); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_243 = 10'hee == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_242); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_244 = 10'hef == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_243); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_245 = 10'hf0 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_244); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_246 = 10'hf1 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_245); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_247 = 10'hf2 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_246); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_248 = 10'hf3 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_247); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_249 = 10'hf4 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_248); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_250 = 10'hf5 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_249); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_251 = 10'hf6 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_250); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_252 = 10'hf7 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_251); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_253 = 10'hf8 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_252); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_254 = 10'hf9 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_253); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_255 = 10'hfa == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_254); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_256 = 10'hfb == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_255); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_257 = 10'hfc == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_256); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_258 = 10'hfd == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_257); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_259 = 10'hfe == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_258); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_260 = 10'hff == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_259); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_261 = 10'h100 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_260); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_262 = 10'h101 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_261); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_263 = 10'h102 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_262); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_264 = 10'h103 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_263); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_265 = 10'h104 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_264); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_266 = 10'h105 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_265); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_267 = 10'h106 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_266); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_268 = 10'h107 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_267); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_269 = 10'h108 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_268); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_270 = 10'h109 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_269); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_271 = 10'h10a == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_270); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_272 = 10'h10b == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_271); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_273 = 10'h10c == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_272); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_274 = 10'h10d == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_273); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_275 = 10'h10e == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_274); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_276 = 10'h10f == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_275); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_277 = 10'h110 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_276); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_278 = 10'h111 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_277); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_279 = 10'h112 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_278); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_280 = 10'h113 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_279); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_281 = 10'h114 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_280); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_282 = 10'h115 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_281); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_283 = 10'h116 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_282); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_284 = 10'h117 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_283); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_285 = 10'h118 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_284); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_286 = 10'h119 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_285); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_287 = 10'h11a == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_286); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_288 = 10'h11b == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_287); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_289 = 10'h11c == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_288); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_290 = 10'h11d == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_289); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_291 = 10'h11e == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_290); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_292 = 10'h11f == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_291); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_293 = 10'h120 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_292); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_294 = 10'h121 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_293); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_295 = 10'h122 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_294); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_296 = 10'h123 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_295); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_297 = 10'h124 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_296); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_298 = 10'h125 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_297); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_299 = 10'h126 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_298); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_300 = 10'h127 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_299); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_301 = 10'h128 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_300); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_302 = 10'h129 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_301); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_303 = 10'h12a == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_302); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_304 = 10'h12b == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_303); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_305 = 10'h12c == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_304); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_306 = 10'h12d == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_305); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_307 = 10'h12e == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_306); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_308 = 10'h12f == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_307); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_309 = 10'h130 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_308); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_310 = 10'h131 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_309); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_311 = 10'h132 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_310); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_312 = 10'h133 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_311); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_313 = 10'h134 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_312); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_314 = 10'h135 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_313); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_315 = 10'h136 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_314); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_316 = 10'h137 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_315); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_317 = 10'h138 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_316); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_318 = 10'h139 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_317); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_319 = 10'h13a == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_318); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_320 = 10'h13b == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_319); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_321 = 10'h13c == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_320); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_322 = 10'h13d == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_321); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_323 = 10'h13e == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_322); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_324 = 10'h13f == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_323); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_325 = 10'h140 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_324); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_326 = 10'h141 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_325); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_327 = 10'h142 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_326); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_328 = 10'h143 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_327); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_329 = 10'h144 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_328); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_330 = 10'h145 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_329); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_331 = 10'h146 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_330); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_332 = 10'h147 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_331); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_333 = 10'h148 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_332); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_334 = 10'h149 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_333); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_335 = 10'h14a == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_334); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_336 = 10'h14b == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_335); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_337 = 10'h14c == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_336); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_338 = 10'h14d == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_337); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_339 = 10'h14e == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_338); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_340 = 10'h14f == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_339); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_341 = 10'h150 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_340); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_342 = 10'h151 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_341); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_343 = 10'h152 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_342); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_344 = 10'h153 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_343); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_345 = 10'h154 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_344); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_346 = 10'h155 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_345); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_347 = 10'h156 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_346); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_348 = 10'h157 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_347); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_349 = 10'h158 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_348); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_350 = 10'h159 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_349); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_351 = 10'h15a == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_350); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_352 = 10'h15b == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_351); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_353 = 10'h15c == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_352); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_354 = 10'h15d == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_353); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_355 = 10'h15e == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_354); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_356 = 10'h15f == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_355); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_357 = 10'h160 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_356); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_358 = 10'h161 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_357); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_359 = 10'h162 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_358); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_360 = 10'h163 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_359); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_361 = 10'h164 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_360); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_362 = 10'h165 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_361); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_363 = 10'h166 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_362); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_364 = 10'h167 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_363); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_365 = 10'h168 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_364); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_366 = 10'h169 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_365); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_367 = 10'h16a == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_366); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_368 = 10'h16b == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_367); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_369 = 10'h16c == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_368); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_370 = 10'h16d == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_369); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_371 = 10'h16e == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_370); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_372 = 10'h16f == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_371); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_373 = 10'h170 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_372); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_374 = 10'h171 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_373); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_375 = 10'h172 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_374); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_376 = 10'h173 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_375); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_377 = 10'h174 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_376); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_378 = 10'h175 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_377); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_379 = 10'h176 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_378); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_380 = 10'h177 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_379); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_381 = 10'h178 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_380); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_382 = 10'h179 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_381); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_383 = 10'h17a == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_382); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_384 = 10'h17b == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_383); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_385 = 10'h17c == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_384); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_386 = 10'h17d == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_385); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_387 = 10'h17e == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_386); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_388 = 10'h17f == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_387); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_389 = 10'h180 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_388); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_390 = 10'h181 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_389); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_391 = 10'h182 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_390); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_392 = 10'h183 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_391); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_393 = 10'h184 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_392); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_394 = 10'h185 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_393); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_395 = 10'h186 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_394); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_396 = 10'h187 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_395); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_397 = 10'h188 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_396); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_398 = 10'h189 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_397); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_399 = 10'h18a == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_398); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_400 = 10'h18b == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_399); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_401 = 10'h18c == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_400); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_402 = 10'h18d == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_401); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_403 = 10'h18e == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_402); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_404 = 10'h18f == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_403); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_405 = 10'h190 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_404); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_406 = 10'h191 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_405); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_407 = 10'h192 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_406); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_408 = 10'h193 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_407); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_409 = 10'h194 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_408); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_410 = 10'h195 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_409); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_411 = 10'h196 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_410); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_412 = 10'h197 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_411); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_413 = 10'h198 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_412); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_414 = 10'h199 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_413); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_415 = 10'h19a == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_414); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_416 = 10'h19b == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_415); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_417 = 10'h19c == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_416); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_418 = 10'h19d == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_417); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_419 = 10'h19e == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_418); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_420 = 10'h19f == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_419); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_421 = 10'h1a0 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_420); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_422 = 10'h1a1 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_421); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_423 = 10'h1a2 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_422); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_424 = 10'h1a3 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_423); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_425 = 10'h1a4 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_424); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_426 = 10'h1a5 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_425); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_427 = 10'h1a6 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_426); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_428 = 10'h1a7 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_427); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_429 = 10'h1a8 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_428); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_430 = 10'h1a9 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_429); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_431 = 10'h1aa == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_430); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_432 = 10'h1ab == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_431); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_433 = 10'h1ac == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_432); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_434 = 10'h1ad == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_433); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_435 = 10'h1ae == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_434); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_436 = 10'h1af == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_435); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_437 = 10'h1b0 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_436); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_438 = 10'h1b1 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_437); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_439 = 10'h1b2 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_438); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_440 = 10'h1b3 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_439); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_441 = 10'h1b4 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_440); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_442 = 10'h1b5 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_441); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_443 = 10'h1b6 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_442); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_444 = 10'h1b7 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_443); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_445 = 10'h1b8 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_444); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_446 = 10'h1b9 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_445); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_447 = 10'h1ba == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_446); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_448 = 10'h1bb == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_447); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_449 = 10'h1bc == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_448); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_450 = 10'h1bd == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_449); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_451 = 10'h1be == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_450); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_452 = 10'h1bf == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_451); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_453 = 10'h1c0 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_452); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_454 = 10'h1c1 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_453); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_455 = 10'h1c2 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_454); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_456 = 10'h1c3 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_455); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_457 = 10'h1c4 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_456); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_458 = 10'h1c5 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_457); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_459 = 10'h1c6 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_458); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_460 = 10'h1c7 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_459); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_461 = 10'h1c8 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_460); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_462 = 10'h1c9 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_461); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_463 = 10'h1ca == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_462); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_464 = 10'h1cb == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_463); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_465 = 10'h1cc == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_464); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_466 = 10'h1cd == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_465); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_467 = 10'h1ce == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_466); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_468 = 10'h1cf == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_467); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_469 = 10'h1d0 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_468); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_470 = 10'h1d1 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_469); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_471 = 10'h1d2 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_470); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_472 = 10'h1d3 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_471); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_473 = 10'h1d4 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_472); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_474 = 10'h1d5 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_473); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_475 = 10'h1d6 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_474); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_476 = 10'h1d7 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_475); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_477 = 10'h1d8 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_476); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_478 = 10'h1d9 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_477); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_479 = 10'h1da == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_478); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_480 = 10'h1db == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_479); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_481 = 10'h1dc == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_480); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_482 = 10'h1dd == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_481); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_483 = 10'h1de == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_482); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_484 = 10'h1df == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_483); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_485 = 10'h1e0 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_484); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_486 = 10'h1e1 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_485); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_487 = 10'h1e2 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_486); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_488 = 10'h1e3 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_487); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_489 = 10'h1e4 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_488); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_490 = 10'h1e5 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_489); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_491 = 10'h1e6 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_490); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_492 = 10'h1e7 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_491); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_493 = 10'h1e8 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_492); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_494 = 10'h1e9 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_493); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_495 = 10'h1ea == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_494); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_496 = 10'h1eb == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_495); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_497 = 10'h1ec == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_496); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_498 = 10'h1ed == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_497); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_499 = 10'h1ee == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_498); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_500 = 10'h1ef == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_499); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_501 = 10'h1f0 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_500); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_502 = 10'h1f1 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_501); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_503 = 10'h1f2 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_502); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_504 = 10'h1f3 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_503); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_505 = 10'h1f4 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_504); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_506 = 10'h1f5 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_505); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_507 = 10'h1f6 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_506); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_508 = 10'h1f7 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_507); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_509 = 10'h1f8 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_508); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_510 = 10'h1f9 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_509); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_511 = 10'h1fa == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_510); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_512 = 10'h1fb == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_511); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_513 = 10'h1fc == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_512); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_514 = 10'h1fd == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_513); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_515 = 10'h1fe == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_514); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_516 = 10'h1ff == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_515); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_517 = 10'h200 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_516); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_518 = 10'h201 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_517); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_519 = 10'h202 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_518); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_520 = 10'h203 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_519); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_521 = 10'h204 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_520); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_522 = 10'h205 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_521); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_523 = 10'h206 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_522); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_524 = 10'h207 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_523); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_525 = 10'h208 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_524); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_526 = 10'h209 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_525); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_527 = 10'h20a == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_526); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_528 = 10'h20b == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_527); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_529 = 10'h20c == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_528); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_530 = 10'h20d == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_529); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_531 = 10'h20e == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_530); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_532 = 10'h20f == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_531); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_533 = 10'h210 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_532); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_534 = 10'h211 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_533); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_535 = 10'h212 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_534); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_536 = 10'h213 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_535); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_537 = 10'h214 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_536); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_538 = 10'h215 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_537); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_539 = 10'h216 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_538); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_540 = 10'h217 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_539); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_541 = 10'h218 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_540); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_542 = 10'h219 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_541); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_543 = 10'h21a == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_542); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_544 = 10'h21b == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_543); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_545 = 10'h21c == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_544); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_546 = 10'h21d == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_545); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_547 = 10'h21e == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_546); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_548 = 10'h21f == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_547); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_549 = 10'h220 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_548); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_550 = 10'h221 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_549); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_551 = 10'h222 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_550); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_552 = 10'h223 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_551); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_553 = 10'h224 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_552); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_554 = 10'h225 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_553); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_555 = 10'h226 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_554); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_556 = 10'h227 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_555); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_557 = 10'h228 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_556); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_558 = 10'h229 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_557); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_559 = 10'h22a == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_558); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_560 = 10'h22b == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_559); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_561 = 10'h22c == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_560); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_562 = 10'h22d == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_561); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_563 = 10'h22e == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_562); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_564 = 10'h22f == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_563); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_565 = 10'h230 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_564); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_566 = 10'h231 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_565); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_567 = 10'h232 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_566); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_568 = 10'h233 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_567); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_569 = 10'h234 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_568); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_570 = 10'h235 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_569); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_571 = 10'h236 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_570); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_572 = 10'h237 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_571); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_573 = 10'h238 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_572); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_574 = 10'h239 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_573); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_575 = 10'h23a == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_574); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_576 = 10'h23b == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_575); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_577 = 10'h23c == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_576); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_578 = 10'h23d == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_577); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_579 = 10'h23e == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_578); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_580 = 10'h23f == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_579); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_581 = 10'h240 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_580); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_582 = 10'h241 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_581); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_583 = 10'h242 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_582); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_584 = 10'h243 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_583); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_585 = 10'h244 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_584); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_586 = 10'h245 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_585); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_587 = 10'h246 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_586); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_588 = 10'h247 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_587); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_589 = 10'h248 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_588); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_590 = 10'h249 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_589); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_591 = 10'h24a == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_590); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_592 = 10'h24b == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_591); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_593 = 10'h24c == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_592); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_594 = 10'h24d == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_593); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_595 = 10'h24e == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_594); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_596 = 10'h24f == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_595); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_597 = 10'h250 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_596); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_598 = 10'h251 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_597); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_599 = 10'h252 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_598); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_600 = 10'h253 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_599); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_601 = 10'h254 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_600); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_602 = 10'h255 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_601); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_603 = 10'h256 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_602); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_604 = 10'h257 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_603); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_605 = 10'h258 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_604); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_606 = 10'h259 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_605); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_607 = 10'h25a == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_606); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_608 = 10'h25b == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_607); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_609 = 10'h25c == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_608); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_610 = 10'h25d == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_609); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_611 = 10'h25e == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_610); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_612 = 10'h25f == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_611); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_613 = 10'h260 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_612); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_614 = 10'h261 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_613); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_615 = 10'h262 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_614); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_616 = 10'h263 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_615); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_617 = 10'h264 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_616); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_618 = 10'h265 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_617); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_619 = 10'h266 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_618); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_620 = 10'h267 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_619); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_621 = 10'h268 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_620); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_622 = 10'h269 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_621); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_623 = 10'h26a == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_622); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_624 = 10'h26b == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_623); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_625 = 10'h26c == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_624); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_626 = 10'h26d == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_625); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_627 = 10'h26e == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_626); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_628 = 10'h26f == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_627); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_629 = 10'h270 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_628); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_630 = 10'h271 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_629); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_631 = 10'h272 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_630); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_632 = 10'h273 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_631); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_633 = 10'h274 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_632); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_634 = 10'h275 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_633); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_635 = 10'h276 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_634); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_636 = 10'h277 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_635); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_637 = 10'h278 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_636); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_638 = 10'h279 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_637); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_639 = 10'h27a == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_638); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_640 = 10'h27b == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_639); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_641 = 10'h27c == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_640); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_642 = 10'h27d == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_641); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_643 = 10'h27e == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_642); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_644 = 10'h27f == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_643); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_645 = 10'h280 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_644); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_646 = 10'h281 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_645); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_647 = 10'h282 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_646); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_648 = 10'h283 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_647); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_649 = 10'h284 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_648); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_650 = 10'h285 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_649); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_651 = 10'h286 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_650); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_652 = 10'h287 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_651); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_653 = 10'h288 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_652); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_654 = 10'h289 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_653); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_655 = 10'h28a == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_654); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_656 = 10'h28b == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_655); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_657 = 10'h28c == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_656); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_658 = 10'h28d == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_657); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_659 = 10'h28e == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_658); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_660 = 10'h28f == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_659); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_661 = 10'h290 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_660); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_662 = 10'h291 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_661); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_663 = 10'h292 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_662); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_664 = 10'h293 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_663); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_665 = 10'h294 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_664); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_666 = 10'h295 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_665); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_667 = 10'h296 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_666); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_668 = 10'h297 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_667); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_669 = 10'h298 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_668); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_670 = 10'h299 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_669); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_671 = 10'h29a == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_670); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_672 = 10'h29b == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_671); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_673 = 10'h29c == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_672); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_674 = 10'h29d == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_673); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_675 = 10'h29e == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_674); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_676 = 10'h29f == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_675); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_677 = 10'h2a0 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_676); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_678 = 10'h2a1 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_677); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_679 = 10'h2a2 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_678); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_680 = 10'h2a3 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_679); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_681 = 10'h2a4 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_680); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_682 = 10'h2a5 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_681); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_683 = 10'h2a6 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_682); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_684 = 10'h2a7 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_683); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_685 = 10'h2a8 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_684); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_686 = 10'h2a9 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_685); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_687 = 10'h2aa == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_686); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_688 = 10'h2ab == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_687); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_689 = 10'h2ac == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_688); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_690 = 10'h2ad == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_689); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_691 = 10'h2ae == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_690); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_692 = 10'h2af == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_691); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_693 = 10'h2b0 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_692); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_694 = 10'h2b1 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_693); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_695 = 10'h2b2 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_694); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_696 = 10'h2b3 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_695); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_697 = 10'h2b4 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_696); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_698 = 10'h2b5 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_697); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_699 = 10'h2b6 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_698); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_700 = 10'h2b7 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_699); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_701 = 10'h2b8 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_700); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_702 = 10'h2b9 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_701); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_703 = 10'h2ba == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_702); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_704 = 10'h2bb == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_703); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_705 = 10'h2bc == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_704); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_706 = 10'h2bd == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_705); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_707 = 10'h2be == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_706); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_708 = 10'h2bf == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_707); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_709 = 10'h2c0 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_708); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_710 = 10'h2c1 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_709); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_711 = 10'h2c2 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_710); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_712 = 10'h2c3 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_711); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_713 = 10'h2c4 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_712); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_714 = 10'h2c5 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_713); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_715 = 10'h2c6 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_714); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_716 = 10'h2c7 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_715); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_717 = 10'h2c8 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_716); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_718 = 10'h2c9 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_717); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_719 = 10'h2ca == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_718); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_720 = 10'h2cb == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_719); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_721 = 10'h2cc == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_720); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_722 = 10'h2cd == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_721); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_723 = 10'h2ce == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_722); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_724 = 10'h2cf == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_723); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_725 = 10'h2d0 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_724); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_726 = 10'h2d1 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_725); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_727 = 10'h2d2 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_726); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_728 = 10'h2d3 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_727); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_729 = 10'h2d4 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_728); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_730 = 10'h2d5 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_729); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_731 = 10'h2d6 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_730); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_732 = 10'h2d7 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_731); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_733 = 10'h2d8 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_732); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_734 = 10'h2d9 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_733); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_735 = 10'h2da == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_734); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_736 = 10'h2db == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_735); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_737 = 10'h2dc == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_736); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_738 = 10'h2dd == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_737); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_739 = 10'h2de == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_738); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_740 = 10'h2df == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_739); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_741 = 10'h2e0 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_740); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_742 = 10'h2e1 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_741); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_743 = 10'h2e2 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_742); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_744 = 10'h2e3 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_743); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_745 = 10'h2e4 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_744); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_746 = 10'h2e5 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_745); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_747 = 10'h2e6 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_746); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_748 = 10'h2e7 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_747); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_749 = 10'h2e8 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_748); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_750 = 10'h2e9 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_749); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_751 = 10'h2ea == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_750); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_752 = 10'h2eb == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_751); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_753 = 10'h2ec == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_752); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_754 = 10'h2ed == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_753); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_755 = 10'h2ee == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_754); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_756 = 10'h2ef == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_755); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_757 = 10'h2f0 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_756); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_758 = 10'h2f1 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_757); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_759 = 10'h2f2 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_758); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_760 = 10'h2f3 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_759); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_761 = 10'h2f4 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_760); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_762 = 10'h2f5 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_761); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_763 = 10'h2f6 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_762); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_764 = 10'h2f7 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_763); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_765 = 10'h2f8 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_764); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_766 = 10'h2f9 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_765); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_767 = 10'h2fa == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_766); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_768 = 10'h2fb == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_767); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_769 = 10'h2fc == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_768); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_770 = 10'h2fd == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_769); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_771 = 10'h2fe == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_770); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_772 = 10'h2ff == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_771); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_773 = 10'h300 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_772); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_774 = 10'h301 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_773); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_775 = 10'h302 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_774); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_776 = 10'h303 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_775); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_777 = 10'h304 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_776); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_778 = 10'h305 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_777); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_779 = 10'h306 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_778); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_780 = 10'h307 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_779); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_781 = 10'h308 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_780); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_782 = 10'h309 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_781); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_783 = 10'h30a == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_782); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_784 = 10'h30b == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_783); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_785 = 10'h30c == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_784); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_786 = 10'h30d == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_785); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_787 = 10'h30e == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_786); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_788 = 10'h30f == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_787); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_789 = 10'h310 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_788); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_790 = 10'h311 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_789); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_791 = 10'h312 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_790); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_792 = 10'h313 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_791); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_793 = 10'h314 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_792); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_794 = 10'h315 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_793); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_795 = 10'h316 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_794); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_796 = 10'h317 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_795); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_797 = 10'h318 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_796); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_798 = 10'h319 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_797); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_799 = 10'h31a == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_798); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_800 = 10'h31b == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_799); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_801 = 10'h31c == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_800); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_802 = 10'h31d == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_801); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_803 = 10'h31e == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_802); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_804 = 10'h31f == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_803); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_805 = 10'h320 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_804); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_806 = 10'h321 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_805); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_807 = 10'h322 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_806); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_808 = 10'h323 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_807); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_809 = 10'h324 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_808); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_810 = 10'h325 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_809); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_811 = 10'h326 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_810); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_812 = 10'h327 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_811); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_813 = 10'h328 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_812); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_814 = 10'h329 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_813); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_815 = 10'h32a == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_814); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_816 = 10'h32b == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_815); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_817 = 10'h32c == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_816); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_818 = 10'h32d == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_817); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_819 = 10'h32e == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_818); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_820 = 10'h32f == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_819); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_821 = 10'h330 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_820); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_822 = 10'h331 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_821); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_823 = 10'h332 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_822); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_824 = 10'h333 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_823); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_825 = 10'h334 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_824); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_826 = 10'h335 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_825); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_827 = 10'h336 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_826); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_828 = 10'h337 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_827); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_829 = 10'h338 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_828); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_830 = 10'h339 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_829); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_831 = 10'h33a == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_830); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_832 = 10'h33b == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_831); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_833 = 10'h33c == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_832); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_834 = 10'h33d == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_833); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_835 = 10'h33e == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_834); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_836 = 10'h33f == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_835); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_837 = 10'h340 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_836); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_838 = 10'h341 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_837); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_839 = 10'h342 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_838); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_840 = 10'h343 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_839); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_841 = 10'h344 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_840); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_842 = 10'h345 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_841); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_843 = 10'h346 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_842); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_844 = 10'h347 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_843); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_845 = 10'h348 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_844); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_846 = 10'h349 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_845); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_847 = 10'h34a == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_846); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_848 = 10'h34b == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_847); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_849 = 10'h34c == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_848); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_850 = 10'h34d == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_849); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_851 = 10'h34e == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_850); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_852 = 10'h34f == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_851); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_853 = 10'h350 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_852); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_854 = 10'h351 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_853); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_855 = 10'h352 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_854); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_856 = 10'h353 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_855); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_857 = 10'h354 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_856); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_858 = 10'h355 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_857); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_859 = 10'h356 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_858); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_860 = 10'h357 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_859); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_861 = 10'h358 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_860); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_862 = 10'h359 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_861); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_863 = 10'h35a == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_862); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_864 = 10'h35b == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_863); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_865 = 10'h35c == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_864); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_866 = 10'h35d == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_865); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_867 = 10'h35e == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_866); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_868 = 10'h35f == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_867); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_869 = 10'h360 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_868); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_870 = 10'h361 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_869); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_871 = 10'h362 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_870); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_872 = 10'h363 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_871); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_873 = 10'h364 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_872); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_874 = 10'h365 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_873); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_875 = 10'h366 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_874); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_876 = 10'h367 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_875); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_877 = 10'h368 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_876); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_878 = 10'h369 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_877); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_879 = 10'h36a == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_878); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_880 = 10'h36b == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_879); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_881 = 10'h36c == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_880); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_882 = 10'h36d == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_881); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_883 = 10'h36e == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_882); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_884 = 10'h36f == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_883); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_885 = 10'h370 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_884); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_886 = 10'h371 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_885); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_887 = 10'h372 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_886); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_888 = 10'h373 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_887); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_889 = 10'h374 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_888); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_890 = 10'h375 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_889); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_891 = 10'h376 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_890); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_892 = 10'h377 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_891); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_893 = 10'h378 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_892); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_894 = 10'h379 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_893); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_895 = 10'h37a == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_894); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_896 = 10'h37b == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_895); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_897 = 10'h37c == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_896); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_898 = 10'h37d == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_897); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_899 = 10'h37e == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_898); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_900 = 10'h37f == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_899); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_901 = 10'h380 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_900); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_902 = 10'h381 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_901); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_903 = 10'h382 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_902); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_904 = 10'h383 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_903); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_905 = 10'h384 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_904); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_906 = 10'h385 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_905); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_907 = 10'h386 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_906); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_908 = 10'h387 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_907); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_909 = 10'h388 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_908); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_910 = 10'h389 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_909); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_911 = 10'h38a == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_910); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_912 = 10'h38b == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_911); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_913 = 10'h38c == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_912); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_914 = 10'h38d == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_913); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_915 = 10'h38e == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_914); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_916 = 10'h38f == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_915); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_917 = 10'h390 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_916); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_918 = 10'h391 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_917); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_919 = 10'h392 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_918); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_920 = 10'h393 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_919); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_921 = 10'h394 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_920); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_922 = 10'h395 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_921); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_923 = 10'h396 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_922); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_924 = 10'h397 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_923); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_925 = 10'h398 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_924); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_926 = 10'h399 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_925); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_927 = 10'h39a == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_926); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_928 = 10'h39b == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_927); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_929 = 10'h39c == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_928); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_930 = 10'h39d == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_929); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_931 = 10'h39e == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_930); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_932 = 10'h39f == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_931); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_933 = 10'h3a0 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_932); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_934 = 10'h3a1 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_933); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_935 = 10'h3a2 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_934); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_936 = 10'h3a3 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_935); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_937 = 10'h3a4 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_936); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_938 = 10'h3a5 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_937); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_939 = 10'h3a6 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_938); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_940 = 10'h3a7 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_939); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_941 = 10'h3a8 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_940); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_942 = 10'h3a9 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_941); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_943 = 10'h3aa == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_942); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_944 = 10'h3ab == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_943); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_945 = 10'h3ac == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_944); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_946 = 10'h3ad == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_945); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_947 = 10'h3ae == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_946); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_948 = 10'h3af == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_947); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_949 = 10'h3b0 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_948); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_950 = 10'h3b1 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_949); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_951 = 10'h3b2 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_950); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_952 = 10'h3b3 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_951); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_953 = 10'h3b4 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_952); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_954 = 10'h3b5 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_953); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_955 = 10'h3b6 == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_954); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_956 = 10'h3b7 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_955); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_957 = 10'h3b8 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_956); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_958 = 10'h3b9 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_957); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_959 = 10'h3ba == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_958); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_960 = 10'h3bb == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_959); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_961 = 10'h3bc == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_960); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_962 = 10'h3bd == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_961); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_963 = 10'h3be == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_962); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_964 = 10'h3bf == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_963); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_965 = 10'h3c0 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_964); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_966 = 10'h3c1 == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_965); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_967 = 10'h3c2 == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_966); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_968 = 10'h3c3 == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_967); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_969 = 10'h3c4 == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_968); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_970 = 10'h3c5 == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_969); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_971 = 10'h3c6 == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_970); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_972 = 10'h3c7 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_971); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_973 = 10'h3c8 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_972); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_974 = 10'h3c9 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_973); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_975 = 10'h3ca == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_974); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_976 = 10'h3cb == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_975); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_977 = 10'h3cc == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_976); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_978 = 10'h3cd == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_977); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_979 = 10'h3ce == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_978); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_980 = 10'h3cf == FRAME_NR[9:0] ? $signed(16'sh0) : $signed(_GEN_979); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_981 = 10'h3d0 == FRAME_NR[9:0] ? $signed(16'sh2e04) : $signed(_GEN_980); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_982 = 10'h3d1 == FRAME_NR[9:0] ? $signed(-16'sh5592) : $signed(_GEN_981); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_983 = 10'h3d2 == FRAME_NR[9:0] ? $signed(16'sh711a) : $signed(_GEN_982); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_984 = 10'h3d3 == FRAME_NR[9:0] ? $signed(-16'sh7cc1) : $signed(_GEN_983); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_985 = 10'h3d4 == FRAME_NR[9:0] ? $signed(16'sh76e2) : $signed(_GEN_984); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_986 = 10'h3d5 == FRAME_NR[9:0] ? $signed(-16'sh6050) : $signed(_GEN_985); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_987 = 10'h3d6 == FRAME_NR[9:0] ? $signed(16'sh3c38) : $signed(_GEN_986); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_988 = 10'h3d7 == FRAME_NR[9:0] ? $signed(-16'shfab) : $signed(_GEN_987); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_989 = 10'h3d8 == FRAME_NR[9:0] ? $signed(-16'sh1f16) : $signed(_GEN_988); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_990 = 10'h3d9 == FRAME_NR[9:0] ? $signed(16'sh4979) : $signed(_GEN_989); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_991 = 10'h3da == FRAME_NR[9:0] ? $signed(-16'sh698a) : $signed(_GEN_990); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_992 = 10'h3db == FRAME_NR[9:0] ? $signed(16'sh7ac9) : $signed(_GEN_991); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_993 = 10'h3dc == FRAME_NR[9:0] ? $signed(-16'sh7ac9) : $signed(_GEN_992); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_994 = 10'h3dd == FRAME_NR[9:0] ? $signed(16'sh698a) : $signed(_GEN_993); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_995 = 10'h3de == FRAME_NR[9:0] ? $signed(-16'sh4979) : $signed(_GEN_994); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_996 = 10'h3df == FRAME_NR[9:0] ? $signed(16'sh1f16) : $signed(_GEN_995); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_997 = 10'h3e0 == FRAME_NR[9:0] ? $signed(16'shfab) : $signed(_GEN_996); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_998 = 10'h3e1 == FRAME_NR[9:0] ? $signed(-16'sh3c38) : $signed(_GEN_997); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_999 = 10'h3e2 == FRAME_NR[9:0] ? $signed(16'sh6050) : $signed(_GEN_998); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_1000 = 10'h3e3 == FRAME_NR[9:0] ? $signed(-16'sh76e2) : $signed(_GEN_999); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_1001 = 10'h3e4 == FRAME_NR[9:0] ? $signed(16'sh7cc1) : $signed(_GEN_1000); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_1002 = 10'h3e5 == FRAME_NR[9:0] ? $signed(-16'sh711a) : $signed(_GEN_1001); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_1003 = 10'h3e6 == FRAME_NR[9:0] ? $signed(16'sh5592) : $signed(_GEN_1002); // @[Hello.scala 138:{45,45}]
  wire [15:0] _GEN_1004 = 10'h3e7 == FRAME_NR[9:0] ? $signed(-16'sh2e04) : $signed(_GEN_1003); // @[Hello.scala 138:{45,45}]
  wire [31:0] _lutOut_T_1 = {$signed(_GEN_1004), 16'h0}; // @[Hello.scala 138:45]
  wire [31:0] _GEN_2047 = {{16{_GEN_1004[15]}},_GEN_1004}; // @[Hello.scala 138:52]
  wire [31:0] _lutOut_T_5 = $signed(_lutOut_T_1) + $signed(_GEN_2047); // @[Hello.scala 138:52]
  wire [7:0] _bDATA_T_3 = _GEN_2046 - Bit_Counter; // @[Hello.scala 139:46]
  wire [31:0] _bDATA_T_4 = $signed(lutOut) >>> _bDATA_T_3; // @[Hello.scala 139:31]
  wire [31:0] _GEN_2005 = Bit_Counter == 8'h0 | Bit_Counter <= _GEN_2046 ? $signed(_lutOut_T_5) : $signed(lutOut); // @[Hello.scala 134:73 138:22 64:30]
  wire  _GEN_2006 = Bit_Counter == 8'h0 | Bit_Counter <= _GEN_2046 ? _bDATA_T_4[0] : bDATA; // @[Hello.scala 134:73 139:21 62:30]
  wire [31:0] _GEN_2007 = Bit_Counter == 8'h0 | Bit_Counter <= _GEN_2046 ? $signed(lutOut) : $signed({{16{DATA[15]}},
    DATA}); // @[Hello.scala 134:73 140:21 63:30]
  wire [31:0] sw_msb_lsb_16_R = {$signed(io_sw), 16'h0}; // @[Hello.scala 145:43]
  wire [31:0] _GEN_2049 = {{16{io_sw[15]}},io_sw}; // @[Hello.scala 147:52]
  wire [31:0] sw_msb_lsb_32 = $signed(_GEN_2049) + $signed(sw_msb_lsb_16_R); // @[Hello.scala 147:52]
  wire [31:0] _bDATA_T_10 = $signed(sw_msb_lsb_32) >>> _bDATA_T_3; // @[Hello.scala 149:38]
  wire [31:0] _GEN_2008 = $signed(io_sw) == 16'sh0 ? $signed(_GEN_2005) : $signed(lutOut); // @[Hello.scala 132:32 64:30]
  wire  _GEN_2009 = $signed(io_sw) == 16'sh0 ? _GEN_2006 : _bDATA_T_10[0]; // @[Hello.scala 132:32 149:21]
  wire [31:0] _GEN_2010 = $signed(io_sw) == 16'sh0 ? $signed(_GEN_2007) : $signed({{16{io_sw[15]}},io_sw}); // @[Hello.scala 132:32 150:21]
  wire [5:0] _T_15 = 6'h20 / 2'h2; // @[Hello.scala 154:40]
  wire [5:0] _T_17 = _T_15 - 6'h1; // @[Hello.scala 154:47]
  wire [7:0] _GEN_2051 = {{2'd0}, _T_17}; // @[Hello.scala 154:29]
  wire  _GEN_2011 = Bit_Counter >= _GEN_2051 | LRClkr; // @[Hello.scala 154:55 155:20 61:30]
  wire  _T_25 = Bit_Counter == _GEN_2046; // @[Hello.scala 157:71]
  wire  _GEN_2012 = Bit_Counter < _GEN_2051 | Bit_Counter == _GEN_2046 ? 1'h0 : _GEN_2011; // @[Hello.scala 157:91 158:20]
  wire [7:0] _Bit_Counter_T_1 = Bit_Counter + 8'h1; // @[Hello.scala 169:40]
  wire [7:0] _GEN_2013 = _T_25 ? 8'h0 : _Bit_Counter_T_1; // @[Hello.scala 162:48 163:25 169:25]
  wire  _GEN_2016 = current_state & _T_25; // @[Hello.scala 112:28 75:15]
  wire [31:0] _GEN_2019 = current_state ? $signed(_GEN_2010) : $signed({{16{DATA[15]}},DATA}); // @[Hello.scala 112:28 63:30]
  wire  _GEN_2022 = ~current_state ? 1'h0 : current_state; // @[Hello.scala 112:28 116:23]
  wire  _GEN_2023 = ~current_state ? 1'h0 : _GEN_2016; // @[Hello.scala 112:28 117:23]
  wire  _GEN_2024 = ~current_state ? 1'h0 : LRClkr; // @[Hello.scala 112:28 118:23 70:15]
  wire  _GEN_2025 = ~current_state ? 1'h0 : BCLKTckr; // @[Hello.scala 112:28 119:23 69:15]
  wire [15:0] _GEN_2026 = ~current_state ? $signed(16'sh0) : $signed(DATA); // @[Hello.scala 112:28 120:23 72:15]
  wire [7:0] _GEN_2028 = ~current_state ? 8'h0 : Bit_Counter; // @[Hello.scala 112:28 122:23 68:15]
  wire  _GEN_2029 = ~current_state | current_state; // @[Hello.scala 112:28 123:25 56:30]
  wire [31:0] _GEN_2032 = ~current_state ? $signed({{16{DATA[15]}},DATA}) : $signed(_GEN_2019); // @[Hello.scala 112:28 63:30]
  wire  _GEN_2034 = Tckr & _GEN_2022; // @[Hello.scala 110:25 76:15]
  wire [31:0] _GEN_2044 = Tckr ? $signed(_GEN_2032) : $signed({{16{DATA[15]}},DATA}); // @[Hello.scala 110:25 63:30]
  wire [31:0] _GEN_2055 = reset ? $signed(32'sh0) : $signed(_GEN_2044); // @[Hello.scala 63:{30,30}]
  clk_wiz_0_clk_wiz pll ( // @[Hello.scala 47:19]
    .MCLK_48K(pll_MCLK_48K),
    .MCLK_44K(pll_MCLK_44K),
    .locked(pll_locked),
    .clk_in1(pll_clk_in1)
  );
  assign io_Ready = Tckr & _GEN_2023; // @[Hello.scala 110:25 75:15]
  assign io_LRCLK = Tckr ? _GEN_2024 : LRClkr; // @[Hello.scala 110:25 70:15]
  assign io_BCLK = Tckr ? _GEN_2025 : BCLKTckr; // @[Hello.scala 110:25 69:15]
  assign io_MCLK = pll_MCLK_44K; // @[Hello.scala 51:11]
  assign io_DATA = Tckr ? $signed(_GEN_2026) : $signed(DATA); // @[Hello.scala 110:25 72:15]
  assign io_bDATA = bDATA; // @[Hello.scala 71:15]
  assign io_State_o = {{1'd0}, _GEN_2034};
  assign io_BitCntr = Tckr ? _GEN_2028 : Bit_Counter; // @[Hello.scala 110:25 68:15]
  assign io_tick = Tckr; // @[Hello.scala 74:15]
  assign io_CLKR = {{8'd0}, ClkCntr}; // @[Hello.scala 73:15]
  assign pll_clk_in1 = clock; // @[Hello.scala 49:18]
  always @(posedge clock) begin
    if (reset) begin // @[Hello.scala 56:30]
      current_state <= 1'h0; // @[Hello.scala 56:30]
    end else if (Tckr) begin // @[Hello.scala 110:25]
      current_state <= _GEN_2029;
    end
    if (reset) begin // @[Hello.scala 57:30]
      Bit_Counter <= 8'h0; // @[Hello.scala 57:30]
    end else if (Tckr) begin // @[Hello.scala 110:25]
      if (~current_state) begin // @[Hello.scala 112:28]
        Bit_Counter <= 8'h0; // @[Hello.scala 121:23]
      end else if (current_state) begin // @[Hello.scala 112:28]
        Bit_Counter <= _GEN_2013;
      end
    end
    if (reset) begin // @[Hello.scala 58:30]
      ClkCntr <= 8'h0; // @[Hello.scala 58:30]
    end else if (_T_1) begin // @[Hello.scala 91:28]
      ClkCntr <= 8'h0; // @[Hello.scala 94:15]
    end else begin
      ClkCntr <= _ClkCntr_T_1; // @[Hello.scala 81:13]
    end
    if (reset) begin // @[Hello.scala 59:30]
      Tckr <= 1'h0; // @[Hello.scala 59:30]
    end else begin
      Tckr <= _T_1;
    end
    BCLKTckr <= reset | _GEN_0; // @[Hello.scala 60:{30,30}]
    if (reset) begin // @[Hello.scala 61:30]
      LRClkr <= 1'h0; // @[Hello.scala 61:30]
    end else if (Tckr) begin // @[Hello.scala 110:25]
      if (!(~current_state)) begin // @[Hello.scala 112:28]
        if (current_state) begin // @[Hello.scala 112:28]
          LRClkr <= _GEN_2012;
        end
      end
    end
    if (reset) begin // @[Hello.scala 62:30]
      bDATA <= 1'h0; // @[Hello.scala 62:30]
    end else if (Tckr) begin // @[Hello.scala 110:25]
      if (!(~current_state)) begin // @[Hello.scala 112:28]
        if (current_state) begin // @[Hello.scala 112:28]
          bDATA <= _GEN_2009;
        end
      end
    end
    DATA <= _GEN_2055[15:0]; // @[Hello.scala 63:{30,30}]
    if (reset) begin // @[Hello.scala 64:30]
      lutOut <= 32'sh0; // @[Hello.scala 64:30]
    end else if (Tckr) begin // @[Hello.scala 110:25]
      if (!(~current_state)) begin // @[Hello.scala 112:28]
        if (current_state) begin // @[Hello.scala 112:28]
          lutOut <= _GEN_2008;
        end
      end
    end
    if (reset) begin // @[Hello.scala 65:30]
      FRAME_NR <= 16'h0; // @[Hello.scala 65:30]
    end else if (FRAME_NR == 16'hac43) begin // @[Hello.scala 105:32]
      FRAME_NR <= 16'h0; // @[Hello.scala 106:16]
    end else if (io_Ready) begin // @[Hello.scala 101:28]
      FRAME_NR <= _FRAME_NR_T_1; // @[Hello.scala 102:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  current_state = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  Bit_Counter = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  ClkCntr = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  Tckr = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  BCLKTckr = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  LRClkr = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bDATA = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  DATA = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  lutOut = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  FRAME_NR = _RAND_9[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
